`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:06:34 03/13/2016 
// Design Name: 
// Module Name:    sigverifier 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sigverifier(
    input clk,
    input rst_b,
    input start,
    output sigvalid,
    output reg finish
    );

//memory interface
reg mem_sel; //0 --- preserve  1 --- add by 1 
reg [9:0] mem_addr;
wire [1049:0] mem_dout;
reg done; //indicate the end

//timer interface
reg cnt1_sel;  //0 --- reset  1 --- start counting
reg [2:0] cnt1;
reg [1:0] cnt2_sel;  //0 --- reset  1 --- start counting   2 --- hold 
reg [5:0] cnt2;

reg load;

reg [0:9799] shift_reg;
reg	shift_sel;

reg [0:4899] tmp_reg;
reg [1:0] tmp_sel;
wire [0:4899] qc_result;

reg [0:4899] sig_reg;
reg add_sel;



reg [1:0] state;
reg [1:0] next_state;

parameter s_start = 2'd0; parameter s_scan = 2'd1;
parameter s_load = 2'd2; parameter s_finish = 2'd3;

always @(posedge clk) begin
 	if (!rst_b) 
 		state <= s_start;
 	else 
 		state <= next_state;
end

always @(*) begin
	 case (state)
	 	s_start: 
	 		if (start)
		 		next_state = s_load;
	 		else
	 			next_state = s_start;
	 	s_scan: 
	 		if (done)
	 			next_state = s_finish;
	 		else if (cnt2 == 49)
	 			next_state = s_load;
	 		else
	 			next_state = s_scan;				
	 	s_load:
	 		if (cnt1 == 4)
	 			next_state = s_scan;
	 		else 
	 			next_state = s_load;
	 	s_finish: 
	 		next_state = s_finish;
	 endcase
 end

 always @(*) begin
 	case (state)
 		s_start: begin
 			cnt1_sel = 0;
 			cnt2_sel = 0;
 			add_sel = 0;
 			done = 0;
 			shift_sel = 0;
 			finish = 0;
 			if (start)
 				mem_sel = 1;
 			else
 				mem_sel = 0;	
 		end		

 		s_scan: begin	
 			cnt1_sel = 0;
 			cnt2_sel = 1;
 			mem_sel = 0;
 			shift_sel = 1; //scan the input signature
 			tmp_sel = 1; //quasi-cyclic
 			if (mem_addr == 980 && cnt2 == 49)
 				done = 1;
 			else if (shift_reg[0]) begin
 				add_sel = 1;				
 			end
 			else begin
 				add_sel = 0;
 			end

 			if (cnt2 == 49)
 				mem_sel = 1;
 			else
 				mem_sel = 0;	
 		end		
 		s_load: begin
 			//5 steps in total,counted by cnt1
 			add_sel = 0;
 			shift_sel = 0;
 			cnt2_sel = 2; //hold cnt2
 			if (cnt1 != 4) begin
 				mem_sel = 1;
 				cnt1_sel = 1;
 				tmp_sel = 2;
 			end	
 			else begin
 				mem_sel = 0;
  				cnt1_sel = 0;
  				tmp_sel = 3;
  			end		
 		end	
 			
 		s_finish: begin
 			finish = 1'd1;
 			cnt1_sel = 0;
 			cnt2_sel = 0;
 			add_sel = 0;
 			mem_sel = 0;
 			done = 0;
 			shift_sel = 0;
 		end	
 	endcase
 end

//cyclic shift register
always @(posedge clk) begin
	if (!rst_b)
		shift_reg <= 9800'b10100000100100000000010000000000000101000000100000000010000010000000100110100000000000100000000100000000000001010000000000011000000101000110000001000000100000000000000100000100000000000000000000100000011100000000000000100000000000000000000000100000010000000000000000000000000000000000000010000000000000000000000000000100001010000000000000001000100011100100000000000010000000100001000100001000000000000100100000100100000100000000000000010000100000001000010000000000000000000000001100000000010000000011000001000000000000000010000000000001000100000010110001000000000000000000000010010000000000100000000000000100000000000000000001100010000111000000100000000000000000001000000010010000000000000100000000000000100100000000000010000000000000100000000000000000011001000010000000000000100011010000001001100000000000101100000000000000000000000010000001001010010000100000000000000100110000000100000000101000000100110000000000000000000010000000010000000000010000001000000000100000001000100000010000001000000000001000100000000101000101100001000000000000000000000001011000011000000001000001001001100001000000000000000000000000001001000010100010000110000101000000000010001000000000000010000001000000000000000000000100000000000000000100001000000000010000000100100000100100000000000110000000000000000000000000000000010000100000010100000000000000000000000100000000001010000000000000000000000000010000001000000000000000000000000000000000000000001100100100000000001001000000000000100000000001000000000000000000100000000000101100100000000000000001000000000000000000010000000000000001100000000001001010000000010001010100000010000000000000101000001000010000110000100000000000000000000000000000000010010000000000000000010010000000010100000000000000000001000110000000010010000000001000000100000000000000010100101000000000000000000001000000101000000000000010000000000000100000001000101000000000001100010000000100000000000000001000000000000001001001000100000000000000000010110010000000000000000100000000000000000100000000000000100010011100001000000000100000000000000100101000100000000100100000000010000000010010000000000010001011000001000000000001000000000100000000000011001100000000010000001000100010000100000010000000000000000000000000000000000000000000101010010000000000001000000100000000010000000101100101000100000000000010000100100000000001100000100000000100000100000110000010000000000001000000000000011100000000000000000000000001000110100001100000000100100000000000100000001000000110100000000000000000000000000000000000010000001000100000001001000101000010000001010000100110000000010000000000001000000100000001000100000000010110000000000000000010000001000001000000000000000010101000000100000101001000000000011100000000100000000000000010000000100000000000001001100010001000000010010000101000110000000100000000000000000000000000100000000000000000001110000000000000000000000000000000001000000000000000010010010010000000001000100001000001000000000000000010000000010000000000000000010000000101000000000000000000000100000010010000000000001000000000010000000000100000000000010010000000000000001000100000010100000000000000000000000000001000001000000000000000000000010000000010000100000000100100000001100000100000000000000100001100010000000000000100000000000000001001000010101010000000000001011000000000100000010000000000000000000000001001000001001000000010000011100000100000000001000000000001000100000000101001000000010100000001000101000010100010100100010001000000000000000001010001000000000000110000010000000000000000010000000000000001000000000001000000001001000000010000000100000000000100000010000000000000000000000010000000000100000000100000000011100100000000000000100010001000001000000000000000000000000000000000001001010100000010000000010000100000100010000000000000000010000111000000000000000000010000000001000000011000010000000001110000000001000000101000000001000000000000001010000000000010000100000001000000000000000011000100000000000000000100000001100010010000000000010000000000000000000010000000000000000101000010010000000000000010000000000000010010010010100000000000000000000100000000000100000000000000000001000000001000000000000001000000000000000000110000110000000000000000011000010000000100000000000000000000100000000001001001010000000001010000000000000000000000000000000000000000000000001100000000000000000001000100110000000000011000001000001000000010000001100000000000000000000000000001000000010010000000000001000010001000001010000000100000000010000000110000000000010000000000001000001100010000000010110000000000000000011001001000111010010000000110001100100000001111001000100100000000000000100000010000001011000010000000010000100000010000000000000010001000000000000100001001000000000100000010000000000010000100000000000001010000000010101000000000000000000010000000000001100000010000001000001000010000000001000100000000000000010000000000010000000000000100000000000001100100100000000000000010011100001000100000001001001000000100000000000000000000000001000001000010000100001110000000000000000000000000000000000001011100010000000100000000001010110000000000000000000000000010100000000000100000010000110000001000000000000001000001001000000000000001000000000100000011000000000000010011000000000100000010100000001001000000000000100010100010000000000001000000001000000100001000101000000000000001001100010000100001000100000000100000100000100000001000010000000100000000000001000100000010000000000000010000000001000000000110100000000000101001000000011000010000000000000000000000000000000001000000000000000000000100010001000000000100000000000000010000000001010000100000000000000000101100100000001000000000010000010000000000010000000010000100000000000000000011010000000000000100010100010000110000000000000011000100000001000000000100000010000000000100010010010010000000000000000011100000000000000000001000000011000000001000000001000000001000000001000000000010000000000000000000000000000000000101110000000000000100000000110100001000010001000010000110000000000000010000001000010000000000010000001000010000110000000000101110000000000000101000001110000000000000000000100000011000000000010000000000000000000000100000001001000000000000000000000000001000000100000001001000000000000000000010000000010001000000000000000000000000000000001000000000000000000000000000000001000100000000100000000000010000000001000000000000000000100010100000000010100000100000101000000000000001010000000000000000010000000100001000000100000000000000000000000010000001001000000000000000000000000100000000000000000000100100000000100000010011010010000100000000000100000000000000000010000000001000001000000010001000001010010000000000000000000000000000000010000000000000000000001001000000000100001000000100000000100000000101000100000001010000000000000000001000000000100000010000000010100101000000010010000000001000000000000000000000010000110000110001000001000001000000000010000000001000000100000010000001010100000000000010000100000000000100010101000001000001000000000100000000000000010000110010000001010001000000000000000000000100001010100110010000000100001000000000011000000000000100010011010000000001000000000000100000000011001001100000000000000000000100000000000110010000010000010000000000000000001000000000000001100001000010000100000000000000000000000000000000010110000000010011000000000000000100000000100000000000101010000000001000010111000000000000000010000000000100100000000000000000110000000001000000000000000001000000100000000000000000001110000100000010000000010000010000000000000000010100101000000110000000000001000000010110000000001000100000001000000011110000001000010000000000000010000110100010000000000000100000000001010010101000000000000010010010000000000000000010000000001000000000001010110001000010001000000000000000100001000000000000000010001000001000001100010000000000000000000010000011110000000010000010000100010000000000001000100100000000110001000110100000101001000000000000100000000000000100010101000100001000000000000001010001100000001010000000000100000000010001100100000011011000010000000000000000000110000100001000000000000010000000001000010100000001000001000000000001000000100000000100011100000010000001101000000010000000010001010001011000100000000010010000000000000001110110000100000000000010000000000001000001000000001101000000000000000100000110000000000000001000000001000000100000000000000001000010010010000000000000010100000100000000000000000010000001000101000001000001000000000000000000101101000000000000100000000000000000000000001000000000000010000110000000000000000100000000000000000010000100001100100000000000000000001000010100000000000010000000000000010000000000000010000000100000000010000100100100101001000000000000000100001000000100000000000000000000011110000100000000000000000000100000001000000000000000000110110001000000000000001001000000000010000010100000000000000000100000001000000000010100000000101001000000000000010010100000000001001001000101100011001000000000000010010000000011110000000000000000100010000001010000000000000000010000000000000000000000000000001001101000010001000100100001010000000000010010100000000000000000000000000100100000000000000110000001101100010000000000001001011100000000000000011001000000000100100000000100001000000010000000100000010000000001000000001001000000100001010000001000000010000000000000001000100100000000100101000000000000000000010000100000110011000001000100001000100011000000000000000000100000001000000010000000110000000001000000000000000000000000000000000010000000000100001001000000000001010000001000000000000011000000000000000000001101001000010100010001100000000001000000010000000100100000010010101000000000000001000100000000010000000000000000000101000000000000000100000011101110000001000110001000000000000001000000010001000000000001000000100000000000000000000100100000000000000000000000000001000001000000010000000101010000000001000100100000000000001000000110000000010000000001010010100011; //load the signature 
	else if (shift_sel)
		shift_reg <= {shift_reg[1:9799],1'b0};
	else
		shift_reg <= shift_reg;	
end

always @(posedge clk) begin
	if (!rst_b)
		tmp_reg <= 4900'd0;
	else if (tmp_sel == 2'd1) // quasi-cyclic shift 1 bit
		tmp_reg <= qc_result;
	else if (tmp_sel == 2'd2) //shift 1050 bit
		tmp_reg <= {tmp_reg[1050:4899],mem_dout};
	else if (tmp_sel == 2'd3) //shift 700 bit
		tmp_reg <= {tmp_reg[700:4899],mem_dout[1049:350]};
	else
		tmp_reg <= tmp_reg;	
end

//GF(2) adder
always @(posedge clk) begin
	if (!rst_b)
		sig_reg <= 4900'b0; 
	else if (add_sel == 1'd1) // add 
		sig_reg <= tmp_reg ^ sig_reg;
	else 
		sig_reg <= sig_reg;					
end

//integer adder
always @(posedge clk) begin
	if (!rst_b)
		mem_addr <= 10'd0;
	else if (mem_sel == 1'd1)
		mem_addr <= mem_addr + 1'd1;
	else
		mem_addr <= mem_addr;		
end

// counter
always @(posedge clk) begin
	if (!cnt1_sel)
		cnt1 <= 6'd0;
	else
		cnt1 <= cnt1 + 1'd1;		
end

always @(posedge clk) begin
	if (cnt2_sel == 0)
		cnt2 <= 6'd0;
	else if(cnt2_sel == 1)
		cnt2 <= (cnt2 == 49) ? 6'd0 : cnt2 + 1'd1;	
	else 
		cnt2 <= cnt2;		
end


assign sigvalid = sig_reg == 4900'b0000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ? 1'b1 : 1'b0;

//memory blocks
mem_top mem_top(
	//input
	.clk(clk),
	.addr(mem_addr),
	//output
	.dout(mem_dout)
    );

genvar gv_i;

//qc shifter array
generate
	for (gv_i = 0; gv_i < 98; gv_i = gv_i + 1) 
	begin: QC
		qc_shifter qc_shifter(
			.input_vector(tmp_reg[gv_i*50:gv_i*50+49]),
			.output_vector(qc_result[gv_i*50:gv_i*50+49])
			);
	end
endgenerate

endmodule
