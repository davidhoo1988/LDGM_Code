library verilog;
use verilog.vl_types.all;
entity sigverifier_tb is
    generic(
        PERIOD          : integer := 10
    );
end sigverifier_tb;
