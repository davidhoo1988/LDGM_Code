library verilog;
use verilog.vl_types.all;
entity vec_generator_tb is
    generic(
        PERIOD          : integer := 10
    );
end vec_generator_tb;
