`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:59:50 04/01/2016 
// Design Name: 
// Module Name:    vec_generator 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: convert matrix index into a sparse vector 
// <140,10,1>
//////////////////////////////////////////////////////////////////////////////////
module vec_generator(
    input clk,
    input rst_b,
    input start,
    input mode,
    input [13:0] idx,
    output reg finish,
    output [0:9799] vector
    );

reg [13:0] lb, ub, lb_buff, ub_buff;
reg [2:0] lb_sel, ub_sel; // 0 --- hold  1 --- add 10  2 --- add 140    3 --- recover the previous   4 --- add 1 OR minus 130  
reg lb_buff_sel, ub_buff_sel;

reg [0:9799] tmp_reg, tmp_buff_reg;
reg [2:0] tmp_sel; // 0 --- hold  1 --- shift_10  2 --- shift_140   3 --- recover the previous 4 --- shift_1
reg tmp_buff_sel;   

//FSM 
reg [2:0] state;
reg [2:0] next_state;

reg found;

parameter init = 3'd0; parameter shift_10 = 3'd1;
parameter shift_140 = 3'd2; parameter shift_1 = 3'd3;


always @(posedge clk) begin
 	if (!rst_b) 
 		state <= init;
 	else 
 		state <= next_state;
end

always @(*) begin
	 case (state)
	 	init: 
	 		if (start && mode == 0)
		 		next_state = shift_10;
	 		else if (start && mode == 1)
	 			next_state = shift_140;
	 		else
	 			next_state = init;

	 	shift_10:
	 		if (found)
	 			next_state = shift_1;
	 		else 
	 			next_state = shift_10;

	 	shift_1: 
	 		if (found)
	 			next_state = init;
	 		else
	 			next_state = shift_1;

	 	shift_140:
	 		if (found)
	 			next_state = shift_10;
	 		else
	 			next_state = shift_140;				
	 endcase
end	 

always @(*) begin
 	case (state)
 		init: begin
 		 	lb_buff_sel = 0;
 		 	ub_buff_sel = 0;
 		 	tmp_sel = 0;
 		 	tmp_buff_sel = 0;
 		 	found = 0;
 			lb_sel = 0;
 			ub_sel = 0;
 			finish = 0;
 		end

 		shift_10: begin
 			if ((lb == idx || lb < idx) && (ub > idx)) begin
 				found = 1;
 				lb_sel = 0;
 				ub_sel = 0;
 				tmp_sel = 0;
 				if (mode == 0) begin // record a copy of the range for mode-0
 					tmp_buff_sel = 1;
 					lb_buff_sel = 1;
 		 			ub_buff_sel = 1;
 		 		end
 		 		else begin
 		 			tmp_buff_sel = 0;
 					lb_buff_sel = 0;
 		 			ub_buff_sel = 0;		 			
 		 		end 		 		
 			end
 				
 			else begin
 				found = 0;	
 				lb_sel = 1;
 				ub_sel = 1;
 				tmp_sel = 1;
 				lb_buff_sel = 0;
 		 		ub_buff_sel = 0;
 		 		tmp_buff_sel = 0;
 			end
 			finish = 0;
 		end

 		shift_1: begin
 			if (lb == idx) begin //the idx found
 				found = 1;
 				lb_sel = 3; //recover the copy
 				ub_sel = 3; //recover
 				tmp_sel = 3; //recover
 				lb_buff_sel = 0;
 				ub_buff_sel = 0;
 				tmp_buff_sel = 0;
 				finish = 1;
 			end
 			else begin
 				found = 0;
 				lb_sel = 4; // +1
 				ub_sel = 0;
 				tmp_sel = 4;
 				lb_buff_sel = 0;
 				ub_buff_sel = 0;
 				tmp_buff_sel = 0;
 				finish = 0;
 			end
 		end

 		shift_140: begin
 			if ((lb == idx || lb < idx) && (ub > idx)) begin //found then go to shift_10
 				found = 1;
 				lb_sel = 0;
 				ub_sel = 4;
 				tmp_sel = 0;
				// we need to record a copy of mode-1
 				tmp_buff_sel = 1;
 				lb_buff_sel = 1;
 				ub_buff_sel = 1;
 				end	
 			else begin
 				found = 0;
 				lb_sel = 2;
 				ub_sel = 2;
 				tmp_sel = 2;
 				tmp_buff_sel = 0;
 				lb_buff_sel = 0;
 				ub_buff_sel = 0;
 			end
 			finish = 0;
 		end

 	endcase
 end				

//tmp_reg generate the vector
always @(posedge clk) begin
	if (!rst_b)
		tmp_reg <= 9800'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	else if (tmp_sel == 3'd1)//shift 10-bit
		tmp_reg <= {10'b0,tmp_reg[0:9789]};		
	else if (tmp_sel == 3'd2)//shift 140-bit
		tmp_reg <= {140'b0,tmp_reg[0:9659]};
	else if (tmp_sel == 3'd3)	
		tmp_reg <= tmp_buff_reg;	
	else if (tmp_sel == 3'd4)
		tmp_reg <= {1'b0,tmp_reg[0:9798]};
	else
		tmp_reg <= tmp_reg;				
end

always @(posedge clk) begin
	if (!rst_b)
		tmp_buff_reg <= 9800'b0;
	else if (tmp_buff_sel)
		tmp_buff_reg <= tmp_reg;
	else
		tmp_buff_reg <= tmp_buff_reg;	
end

//lower bound reg
always @(posedge clk) begin
	if (!rst_b)
		lb <= 0;
	else if (lb_sel == 3'd1) 
		lb <= lb + 10;
	else if (lb_sel == 3'd2)  
		lb <= lb + 140;
	else if (lb_sel == 3'd3) 
		lb <= lb_buff;	
	else if (lb_sel == 3'd4)
		lb <= lb + 1;	
	else
		lb <= lb;			
end

always @(posedge clk) begin
	if (!rst_b)
		lb_buff <= 0;
	else if (lb_buff_sel)
		lb_buff <= lb; 	
	else
		lb_buff <= lb_buff;
end

//upper bound reg
always @(posedge clk) begin
	if (!rst_b && mode==0)
		ub <= 10;
	else if (!rst_b && mode==1)
		ub <= 140;	
	else if (ub_sel == 3'd1)
		ub <= ub + 10;
	else if (ub_sel == 3'd2) 
		ub <= ub + 140;	
	else if (ub_sel == 3'd3)
		ub <= ub_buff;	
	else if (ub_sel == 3'd4) 
		ub <= ub - 130;
	else
		ub <= ub;	
end

always @(posedge clk) begin
	if (!rst_b)
		ub_buff <= 0;
	else if (ub_buff_sel)
		ub_buff <= ub; 	
	else
		ub_buff <= ub_buff;
end

assign vector = tmp_reg;
endmodule
